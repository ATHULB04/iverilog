module hello();

initial
  begin
    $display("Hello World!");   // This will display a message
  end

endmodule