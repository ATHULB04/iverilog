module sample(a,b,e);
input a,b;
output e;
and a1(e,a,b);
endmodule
